LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY Sub_Bytes_ROM IS
    PORT (
        clock : IN STD_LOGIC;
        address : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
        data_out : OUT STD_LOGIC_VECTOR(8 DOWNTO 0));
END ENTITY;

ARCHITECTURE Sub_Bytes_ROM_ARC OF Sub_Bytes_ROM IS

    TYPE ROM_type IS ARRAY(0 TO 255) OF STD_LOGIC_VECTOR(7 DOWNTO 0);

    CONSTANT ROM : ROM_type := (
        1 => x"63",
        2 => x"7c",
        3 => x"77",
        4 => x"7b",
        5 => x"f2",
        6 => x"6b",
        7 => x"6f",
        8 => x"c5",
        9 => x"30",
        10 => x"01",
        11 => x"67",
        12 => x"2b",
        13 => x"fe",
        14 => x"d7",
        15 => x"ab",
        16 => x"76",
        17 => x"ca",
        18 => x"82",
        19 => x"c9",
        20 => x"7d",
        21 => x"fa",
        22 => x"59",
        23 => x"47",
        24 => x"f0",
        25 => x"ad",
        26 => x"d4",
        27 => x"a2",
        28 => x"af",
        29 => x"9c",
        30 => x"a4",
        31 => x"72",
        32 => x"c0",
        33 => x"b7",
        34 => x"fd",
        35 => x"93",
        36 => x"26",
        37 => x"36",
        38 => x"3f",
        39 => x"f7",
        40 => x"cc",
        41 => x"34",
        42 => x"a5",
        43 => x"e5",
        44 => x"f1",
        45 => x"71",
        46 => x"d8",
        47 => x"31",
        48 => x"15",
        49 => x"04",
        50 => x"c7",
        51 => x"23",
        52 => x"c3",
        53 => x"18",
        54 => x"96",
        55 => x"05",
        56 => x"9a",
        57 => x"07",
        58 => x"12",
        59 => x"80",
        60 => x"e2",
        61 => x"eb",
        62 => x"27",
        63 => x"b2",
        64 => x"75",
        65 => x"09",
        66 => x"83",
        67 => x"2c",
        68 => x"1a",
        69 => x"1b",
        70 => x"6e",
        71 => x"5a",
        72 => x"a0",
        73 => x"52",
        74 => x"3b",
        75 => x"d6",
        76 => x"b3",
        77 => x"29",
        78 => x"e3",
        79 => x"2f",
        80 => x"84",
        81 => x"53",
        82 => x"d1",
        83 => x"00",
        84 => x"ed",
        85 => x"20",
        86 => x"fc",
        87 => x"b1",
        88 => x"5b",
        89 => x"6a",
        90 => x"cb",
        91 => x"be",
        92 => x"39",
        93 => x"4a",
        94 => x"4c",
        95 => x"58",
        96 => x"cf",
        97 => x"d0",
        98 => x"ef",
        99 => x"aa",
        100 => x"fb",
        101 => x"43",
        102 => x"4d",
        103 => x"33",
        104 => x"85",
        105 => x"45",
        106 => x"f9",
        107 => x"02",
        108 => x"7f",
        109 => x"50",
        110 => x"3c",
        111 => x"9f",
        112 => x"a8",
        113 => x"51",
        114 => x"a3",
        115 => x"40",
        116 => x"8f",
        117 => x"92",
        118 => x"9d",
        119 => x"38",
        120 => x"f5",
        121 => x"bc",
        122 => x"b6",
        123 => x"da",
        124 => x"21",
        125 => x"10",
        126 => x"ff",
        127 => x"f3",
        128 => x"d2",
        129 => x"cd",
        130 => x"0c",
        131 => x"13",
        132 => x"ec",
        133 => x"5f",
        134 => x"97",
        135 => x"44",
        136 => x"17",
        137 => x"c4",
        138 => x"a7",
        139 => x"7e",
        140 => x"3d",
        141 => x"64",
        142 => x"5d",
        143 => x"19",
        144 => x"73",
        145 => x"60",
        146 => x"81",
        147 => x"4f",
        148 => x"dc",
        149 => x"22",
        150 => x"2a",
        151 => x"90",
        152 => x"88",
        153 => x"46",
        154 => x"ee",
        155 => x"b8",
        156 => x"14",
        157 => x"de",
        158 => x"5e",
        159 => x"0b",
        160 => x"db",
        161 => x"e0",
        162 => x"32",
        163 => x"3a",
        164 => x"0a",
        165 => x"49",
        166 => x"06",
        167 => x"24",
        168 => x"5c",
        169 => x"c2",
        170 => x"d3",
        171 => x"ac",
        172 => x"62",
        173 => x"91",
        174 => x"95",
        175 => x"e4",
        176 => x"79",
        177 => x"e7",
        178 => x"c8",
        179 => x"37",
        180 => x"6d",
        181 => x"8d",
        182 => x"d5",
        183 => x"4e",
        184 => x"a9",
        185 => x"6c",
        186 => x"56",
        187 => x"f4",
        188 => x"ea",
        189 => x"65",
        190 => x"7a",
        191 => x"ae",
        192 => x"08",
        193 => x"ba",
        194 => x"78",
        195 => x"25",
        196 => x"2e",
        197 => x"1c",
        198 => x"a6",
        199 => x"b4",
        200 => x"c6",
        201 => x"e8",
        202 => x"dd",
        203 => x"74",
        204 => x"1f",
        205 => x"4b",
        206 => x"bd",
        207 => x"8b",
        208 => x"8a",
        209 => x"70",
        210 => x"3e",
        211 => x"b5",
        212 => x"66",
        213 => x"48",
        214 => x"03",
        215 => x"f6",
        216 => x"0e",
        217 => x"61",
        218 => x"35",
        219 => x"57",
        220 => x"b9",
        221 => x"86",
        222 => x"c1",
        223 => x"1d",
        224 => x"9e",
        225 => x"e1",
        226 => x"f8",
        227 => x"98",
        228 => x"11",
        229 => x"69",
        230 => x"d9",
        231 => x"8e",
        232 => x"94",
        233 => x"9b",
        234 => x"1e",
        235 => x"87",
        236 => x"e9",
        237 => x"ce",
        238 => x"55",
        239 => x"28",
        240 => x"df",
        241 => x"8c",
        242 => x"a1",
        243 => x"89",
        244 => x"0d",
        245 => x"bf",
        246 => x"e6",
        247 => x"42",
        248 => x"68",
        249 => x"41",
        250 => x"99",
        251 => x"2d",
        252 => x"0f",
        253 => x"b0",
        254 => x"54",
        255 => x"bb",
        256 => x"16");

BEGIN

    MEMORY : PROCESS (clock)
    BEGIN
        IF (rising_edge(clock)) THEN
            data_out <= ROM(to_integer(unsigned(address)));
        END IF;
    END PROCESS;
END ARCHITECTURE;